`timescale 1ns / 1ps

package package_gpr_destination_selector;
  typedef enum logic [3:0] {
    GPR_DESTINATION_SELECTOR_GPR0 = 4'b0000,
    GPR_DESTINATION_SELECTOR_GPR1 = 4'b0001,
    GPR_DESTINATION_SELECTOR_GPR2 = 4'b0010,
    GPR_DESTINATION_SELECTOR_GPR3 = 4'b0011,
    GPR_DESTINATION_SELECTOR_GPR4 = 4'b0100,
    GPR_DESTINATION_SELECTOR_GPR5 = 4'b0101,
    GPR_DESTINATION_SELECTOR_GPR6 = 4'b0110,
    GPR_DESTINATION_SELECTOR_GPR7 = 4'b0111,
    GPR_DESTINATION_SELECTOR_RA   = 4'b1000,
    GPR_DESTINATION_SELECTOR_RAP  = 4'b1001,
    GPR_DESTINATION_SELECTOR_RB   = 4'b1010,
    GPR_DESTINATION_SELECTOR_RBP  = 4'b1011,
    GPR_DESTINATION_SELECTOR_NONE = 4'b1111
  } GPR_DESTINATION_SELECTOR;
endpackage
