`timescale 1ns / 1ps

package package_control_data;
  typedef logic [39:0] MICRO1_CONTROL_WORD;
  typedef logic [11:0] MICRO1_CONTROL_ADDRESS;
endpackage
