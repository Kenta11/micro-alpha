`timescale 1ns / 1ps

package package_machine_data;
  typedef logic [15:0] MICRO1_MACHINE_WORD;
  typedef logic [15:0] MICRO1_MACHINE_ADDRESS;
endpackage
